//axi write related
`define AXI_OKAY                    2'b00
`define AXI_EXOKAY                  2'b01
`define AXI_SLVERR                  2'b10
`define AXI_DECERR                  2'b11
// burst type
`define AXI_WR_BURST_FIXED          2'b00
`define AXI_WR_BURST_INCR           2'b01
`define AXI_WR_BURST_WRAP           2'b10
// region define
`define AXI_CMD_FIFO_REGION         4'b0
`define AXI_WRAM_REGION             4'b1
`define AXI_IRAM_REGION             4'b10
// max values
`define AWBURST_MAX                 3'b010

`define CMD_MSB                     63
`define CMD_OP_WIDTH                5
`define CMD_OP_LSB                  (CMD_MSB-CMD_OP_WIDTH+1)

`define CMD_WRAM_ADDR_WIDTH         8
`define CMD_WRAM_ADDR_MSB           (CMD_OP_LSB-1)
`define CMD_WRAM_ADDR_LSB           (CMD_WRAM_ADDR_MSB-CMD_WRAM_ADDR_WIDTH+1)
`define CMD_WRAM_ADDR_RNG           CMD_WRAM_ADDR_MSB:CMD_WRAM_ADDR_LSB

`define CMD_WRAM_START_ADDR_WIDTH   4
`define CMD_WRAM_START_ADDR_MSB     (CMD_WRAM_ADDR_LSB-1)
`define CMD_WRAM_START_ADDR_LSB     (CMD_WRAM_START_ADDR_MSB-CMD_WRAM_START_ADDR_WIDTH+1)
`define CMD_WRAM_START_ADDR_RNG     CMD_WRAM_START_ADDR_MSB:CMD_WRAM_START_ADDR_LSB

`define CMD_WRAM_END_ADDR_WIDTH     4
`define CMD_WRAM_END_ADDR_MSB       (CMD_WRAM_START_ADDR_LSB-1)
`define CMD_WRAM_END_ADDR_LSB       (CMD_WRAM_END_ADDR_MSB-CMD_WRAM_END_ADDR_WIDTH+1)
`define CMD_WRAM_END_ADDR_RNG       CMD_WRAM_END_ADDR_MSB:CMD_WRAM_END_ADDR_LSB

`define CMD_IRAM_ADDR_WIDTH         8
`define CMD_IRAM_ADDR_MSB           (CMD_WRAM_END_ADDR_LSB-1)
`define CMD_IRAM_ADDR_LSB           (CMD_IRAM_ADDR_MSB-CMD_IRAM_ADDR_WIDTH+1)
`define CMD_IRAM_ADDR_RNG           CMD_IRAM_ADDR_MSB:CMD_IRAM_ADDR_LSB

`define CMD_IRAM_START_ADDR_WIDTH   4
`define CMD_IRAM_START_ADDR_MSB     (CMD_IRAM_ADDR_LSB-1)
`define CMD_IRAM_START_ADDR_LSB     (CMD_IRAM_START_ADDR_MSB-CMD_IRAM_START_ADDR_WIDTH+1)
`define CMD_IRAM_START_ADDR_RNG     CMD_IRAM_START_ADDR_MSB:CMD_IRAM_START_ADDR_LSB

`define CMD_IRAM_END_ADDR_WIDTH     4
`define CMD_IRAM_END_ADDR_MSB       (CMD_IRAM_START_ADDR_LSB-1)
`define CMD_IRAM_END_ADDR_LSB       (CMD_IRAM_END_ADDR_MSB-CMD_IRAM_END_ADDR_WIDTH+1)
`define CMD_IRAM_END_ADDR_RNG       CMD_IRAM_END_ADDR_MSB:CMD_IRAM_END_ADDR_LSB

`define CMD_ORAM_ADDR_WIDTH         8
`define CMD_ORAM_ADDR_MSB           (CMD_IRAM_END_ADDR_LSB-1)
`define CMD_ORAM_ADDR_LSB           (CMD_ORAM_ADDR_MSB-CMD_ORAM_ADDR_WIDTH+1)
`define CMD_ORAM_ADDR_RNG           CMD_ORAM_ADDR_MSB:CMD_ORAM_ADDR_LSB

`define CMD_ORAM_START_ADDR_WIDTH   4
`define CMD_ORAM_START_ADDR_MSB     (CMD_ORAM_ADDR_LSB-1)
`define CMD_ORAM_START_ADDR_LSB     (CMD_ORAM_START_ADDR_MSB-CMD_ORAM_START_ADDR_WIDTH+1)
`define CMD_ORAM_START_ADDR_RNG     CMD_ORAM_START_ADDR_MSB:CMD_ORAM_START_ADDR_LSB

`define CMD_ORAM_END_ADDR_WIDTH     4
`define CMD_ORAM_END_ADDR_MSB       (CMD_ORAM_START_ADDR_LSB-1)
`define CMD_ORAM_END_ADDR_LSB       (CMD_ORAM_END_ADDR_MSB-CMD_ORAM_END_ADDR_WIDTH+1)
`define CMD_ORAM_END_ADDR_RNG       CMD_ORAM_END_ADDR_MSB:CMD_ORAM_END_ADDR_LSB

//RAM buff fsm
`define RAM_BUFF_FSM_IDLE           00
`define RAM_BUFF_FSM_RECV           01
`define RAM_BUFF_FSM_SND            10
`define RAM_BUFF_FSM_REV            11